library verilog;
use verilog.vl_types.all;
entity Mux4_16_vlg_vec_tst is
end Mux4_16_vlg_vec_tst;
